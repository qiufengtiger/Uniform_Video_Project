module tracking_module(
	input clk,
	output azResult,
	output elResult
    );

	assign azResult = 1;
	assign elResult = 1;

endmodule
