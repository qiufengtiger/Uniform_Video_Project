module crosshair_module(
	input vsync,
	input csync,
	input clk4mhz,
	input en,
	input xCounterEn,
	output isCrosshair,
	output [8 : 0] lineCount,
	output [8 : 0] columnCount
    );

	// wire en;
	// wire xCounterEn;


	
	//x & y index
	

	


endmodule
