module cpld_toplevel(
	input vsync,
	input burst,
	input field,
	input csync,
	output gate_b,
	output gate_w
	);


endmodule
